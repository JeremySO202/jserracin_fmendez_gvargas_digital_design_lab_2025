module Sec_conx(
	input logic clk, rst, rx, rx_e, tick,
	input logic[2:0] recep,
	output logic rxReady,
	output logic [7:0] rxOut

);


//2 estados, no leer y leer

parameter IDLE = 1'b0, READ = 1'b1;

reg [1:0] State, Next;

//variables para la maquina

reg read_enable = 1'b0;
reg start_bit = 1'b1;
reg [4:0] Bit = 5'b00000;
reg [3:0] counter = 4'b0000;
reg [7:0] read_data = 8'b00000000;


//primero hay q ver lo que pasa con el leer y no leer
always_ff @(posedge clk or negedge rst) begin
	if (!rst)
    State <= IDLE;
	else
    State <= Next;
end

always_comb begin
	case (State)
		IDLE:  Next = (!rx && rx_e) ? READ : IDLE;
      READ:  Next = rxReady ? IDLE : READ;
      default: Next = IDLE;
	endcase
end
	 
always_comb begin 
	case(State)
		READ: read_enable = 1'b1;
		IDLE: read_enable = 1'b0;
		default: read_enable = 1'b0;
	endcase
end

//ahora para lo que se recibe

always_ff @(posedge tick) begin
	if (read_enable) begin
		rxReady <= 1'b0;
		counter <= counter + 1;

		//bit de inicio
		if ((counter == 4'd8) && start_bit) begin
			start_bit <= 1'b0;
			counter <= 4'd0;
		end

		// leer
		if ((counter == 4'd15) && !start_bit && (Bit < recep)) begin
			Bit <= Bit + 1;
			read_data <= {rx, read_data[7:1]};
			counter <= 4'd0;
		end

   // ultimo flanco
	if ((counter == 4'd15) && (Bit == recep) && rx) begin
		Bit <= 5'd0;
		rxReady <= 1'b1;
		counter <= 4'd0;
		start_bit <= 1'b1;
		end
	end
end //end del amways com

// la salida
    always_ff @(posedge clk) begin
        case (recep)
            4'd8: rxOut <= read_data;
            4'd7: rxOut <= {1'b0, read_data[7:1]};
            4'd6: rxOut <= {2'b00, read_data[7:2]};
            default: rxOut <= 8'd0;
        endcase
    end

endmodule