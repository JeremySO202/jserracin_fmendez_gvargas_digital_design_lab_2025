module adder ( 
	);
	
	
	
	

endmodule

